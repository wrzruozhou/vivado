`timescale 1ns / 1ps
//****************************************VSCODE PLUG-IN**********************************//
//----------------------------------------------------------------------------------------
// IDE :                   VSCODE     
// VSCODE plug-in version: Verilog-Hdl-Format-2.6.20240622
// VSCODE plug-in author : Jiang Percy
//----------------------------------------------------------------------------------------
//****************************************Copyright (c)***********************************//
// Copyright(C)            WRZ
// All rights reserved     
// File name:              
// Last modified Date:     2024/07/04 18:11:37
// Last Version:           V1.0
// Descriptions:           
//----------------------------------------------------------------------------------------
// Created by:             WRZ
// Created date:           2024/07/04 18:11:37
// mail      :             2350808537@qq.com
// Version:                V1.0
// TEXT NAME:              and_gate.v
// PATH:                   G:\_FPGA\1\rtl\and_gate.v
// Descriptions:           
//                         
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module and_gate(
    input                               A                        ,
    input                               B                        ,

    output                              Y                          
);

//assign相当于一条线，输入A与输入B想与后连接输出Y
    assign                              Y                         = A & B;
                                                                   
                                                                   
endmodule
